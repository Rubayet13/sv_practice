To make the code more simple and readable. 
consider the following example without enumeration. 


enum {RED,YELLOW, GREEN} light_1; 
enum bit [1:0] 