// double forward slash for single line comment 

/* slash and a asterisk for a multiple line comment 
but for to end a multiple line comment 
//i also have to use another * and a forward slash following that will end the multiple line comments
*/


/* there are 4 states basically, 
0,1,x,z
x means it could be either 1 or 0
z means the net has high impedence- maybe the wire is not connected and is floating. 
*/

